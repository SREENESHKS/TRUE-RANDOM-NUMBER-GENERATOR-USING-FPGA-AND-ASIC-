module xor_tree (
    input [31:0] ro_signals,
    output xor_out
);
    assign xor_out = ^ro_signals; // XOR reduction
endmodule
